module teste(input a, input b);
    assign b = a;
endmodule